-- Code your testbench here
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY test_bench IS
END test_bench;

ARCHITECTURE tb_arch OF test_bench IS

    SIGNAL

BEGIN
    mux : ENTITY work.() PORT MAP(
            
        );

    tb_proc : PROCESS

    BEGIN

    END PROCESS;
END tb_arch; -- test_bench